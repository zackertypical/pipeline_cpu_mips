`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:04:38 11/25/2018
// Design Name:   ADD4
// Module Name:   C:/hdl/p5/testadd.v
// Project Name:  p5
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ADD4
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testadd;

	reg  [1:0]in;
	reg [1:0]out;
	reg [1:0]t;
	initial begin
		 out = 0;
		 in = 2;
		 t = 12;//1100
		
		

	end
      
endmodule

